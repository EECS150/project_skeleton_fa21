module bpm_detector();
    // TODO
endmodule
