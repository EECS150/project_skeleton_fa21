module mic_interface();
    // TODO
endmodule
